`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    03:14:31 12/04/2024 
// Design Name: 
// Module Name:    IDO_BUFFER 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module IDO_BUFFER(
    input [15:0] IN_DATA,
    output [15:0] OUT_DATA
    );

assign O = I;


endmodule
