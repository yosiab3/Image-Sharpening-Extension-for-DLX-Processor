`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:53:49 12/08/2024 
// Design Name: 
// Module Name:    BUFFER2BITS 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module BUFFER2BITS(
    input [1:0] IN_D,
    output [1:0] OUT_D
    );

   assign OUT_D = IN_D;


endmodule