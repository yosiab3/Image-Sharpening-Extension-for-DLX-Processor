`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    03:41:17 12/04/2024 
// Design Name: 
// Module Name:    BUFFER_5_BITS 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module BUFFER_5_BITS(
    input [4:0] IN_D,
    output [4:0] OUT_D
    );

   assign OUT_D = IN_D;


endmodule
