`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    03:21:51 12/04/2024 
// Design Name: 
// Module Name:    buffer_4_bytes 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module buffer_4_bytes(
    input [15:0] IN_D,
    output [15:0] OUT_D
    );

   assign OUT_D = IN_D;


endmodule
